module bcd_adder16(a, b, cin, cout, sum);
  input [15:0] a, b;
  input cin;
  output cout;
  output [15:0] sum;
  wire [15:0] a, b;
  wire cin;
  wire cout;
  wire [15:0] sum;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15;
  wire n_16, n_18, n_19, n_20, n_21, n_22, n_23, n_24;
  wire n_25, n_26, n_27, n_29, n_30, n_32, n_33, n_35;
  wire n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44;
  wire n_45, n_46, n_47, n_48, n_50, n_51, n_54, n_56;
  wire n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64;
  wire n_65, n_66, n_67, n_69, n_70, n_73, n_75, n_76;
  wire n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_86;
  wire n_87, n_89, n_90;
  OAI2BB2XL g1161(.A0N (n_89), .A1N (n_90), .B0 (n_90), .B1 (n_89), .Y(sum[15]));
  OAI2BB2XL g1160(.A0N (n_86), .A1N (n_87), .B0 (n_87), .B1 (n_86), .Y(sum[14]));
  OAI21XL g1162(.A0 (cout), .A1 (n_83), .B0 (n_87), .Y (sum[13]));
  NAND2BXL g1163(.AN (n_82), .B (cout), .Y (n_90));
  NAND2XL g1164(.A (n_83), .B (cout), .Y (n_87));
  OAI221XL g1165(.A0 (n_81), .A1 (n_82), .B0 (n_78), .B1 (n_1), .C0(n_0), .Y (cout));
  INVXL g1166(.A (n_89), .Y (n_81));
  OAI2BB2XL g1167(.A0N (n_79), .A1N (n_80), .B0 (n_80), .B1 (n_79), .Y(n_89));
  NOR2XL g1168(.A (n_86), .B (n_76), .Y (n_82));
  OAI21XL g1169(.A0 (n_77), .A1 (n_78), .B0 (n_12), .Y (n_80));
  MXI2XL g1170(.S0 (n_13), .B (n_77), .A (n_75), .Y (n_86));
  INVXL g1171(.A (n_76), .Y (n_83));
  INVXL g1172(.A (n_75), .Y (n_77));
  ADDFX2 g1173(.A (b[13]), .B (a[13]), .CI (n_73), .S (n_76), .CO(n_75));
  ADDFX2 g1176(.A (b[12]), .B (a[12]), .CI (n_62), .S (sum[12]), .CO(n_73));
  DLY4X1 g1175(.A (n_65), .Y (sum[9]));
  OAI2BB2XL g1177(.A0N (n_69), .A1N (n_70), .B0 (n_70), .B1 (n_69), .Y(sum[11]));
  OAI2BB2XL g1174(.A0N (n_66), .A1N (n_67), .B0 (n_67), .B1 (n_66), .Y(sum[10]));
  AOI21XL g1178(.A0 (n_64), .A1 (n_63), .B0 (n_67), .Y (n_65));
  NOR2XL g1179(.A (n_64), .B (n_61), .Y (n_70));
  NOR2XL g1180(.A (n_64), .B (n_63), .Y (n_67));
  INVXL g1181(.A (n_62), .Y (n_64));
  OAI221XL g1182(.A0 (n_69), .A1 (n_61), .B0 (n_58), .B1 (n_3), .C0(n_2), .Y (n_62));
  AOI2BB2XL g1183(.A0N (n_60), .A1N (n_59), .B0 (n_60), .B1 (n_59), .Y(n_69));
  NOR2BXL g1184(.AN (n_66), .B (n_63), .Y (n_61));
  OAI21XL g1185(.A0 (n_57), .A1 (n_58), .B0 (n_10), .Y (n_60));
  MXI2XL g1186(.S0 (n_11), .B (n_56), .A (n_57), .Y (n_66));
  INVXL g1187(.A (n_56), .Y (n_57));
  ADDFX2 g1188(.A (b[9]), .B (a[9]), .CI (n_54), .S (n_63), .CO (n_56));
  ADDFX2 g1191(.A (b[8]), .B (a[8]), .CI (n_43), .S (sum[8]), .CO(n_54));
  INVXL g1190(.A (n_46), .Y (sum[5]));
  OAI2BB2XL g1192(.A0N (n_50), .A1N (n_51), .B0 (n_51), .B1 (n_50), .Y(sum[7]));
  OAI2BB2XL g1189(.A0N (n_47), .A1N (n_48), .B0 (n_48), .B1 (n_47), .Y(sum[6]));
  AOI21XL g1193(.A0 (n_45), .A1 (n_44), .B0 (n_48), .Y (n_46));
  NOR2XL g1194(.A (n_45), .B (n_42), .Y (n_51));
  NOR2XL g1195(.A (n_45), .B (n_44), .Y (n_48));
  INVXL g1196(.A (n_43), .Y (n_45));
  OAI221XL g1197(.A0 (n_50), .A1 (n_42), .B0 (n_39), .B1 (n_9), .C0(n_8), .Y (n_43));
  AOI2BB2XL g1198(.A0N (n_41), .A1N (n_40), .B0 (n_41), .B1 (n_40), .Y(n_50));
  NOR2BXL g1199(.AN (n_47), .B (n_44), .Y (n_42));
  OAI21XL g1200(.A0 (n_38), .A1 (n_39), .B0 (n_14), .Y (n_41));
  MXI2XL g1201(.S0 (n_15), .B (n_37), .A (n_38), .Y (n_47));
  INVXL g1202(.A (n_37), .Y (n_38));
  ADDFX2 g1203(.A (b[5]), .B (a[5]), .CI (n_35), .S (n_44), .CO (n_37));
  ADDFX2 g1206(.A (b[4]), .B (a[4]), .CI (n_24), .S (sum[4]), .CO(n_35));
  OAI2BB2XL g1207(.A0N (n_32), .A1N (n_33), .B0 (n_33), .B1 (n_32), .Y(sum[3]));
  OAI2BB2XL g1204(.A0N (n_29), .A1N (n_30), .B0 (n_30), .B1 (n_29), .Y(sum[2]));
  INVXL g1205(.A (n_27), .Y (sum[1]));
  AOI21XL g1208(.A0 (n_26), .A1 (n_25), .B0 (n_30), .Y (n_27));
  NOR2XL g1209(.A (n_26), .B (n_23), .Y (n_33));
  NOR2XL g1210(.A (n_26), .B (n_25), .Y (n_30));
  INVXL g1211(.A (n_24), .Y (n_26));
  OAI221XL g1212(.A0 (n_32), .A1 (n_23), .B0 (n_19), .B1 (n_5), .C0(n_4), .Y (n_24));
  AOI2BB2XL g1213(.A0N (n_22), .A1N (n_21), .B0 (n_22), .B1 (n_21), .Y(n_32));
  NOR2BXL g1214(.AN (n_29), .B (n_25), .Y (n_23));
  MXI2XL g1216(.S0 (n_7), .B (n_18), .A (n_20), .Y (n_29));
  OAI21XL g1215(.A0 (n_20), .A1 (n_19), .B0 (n_6), .Y (n_22));
  INVXL g1217(.A (n_18), .Y (n_20));
  ADDFX2 g1218(.A (b[1]), .B (a[1]), .CI (n_16), .S (n_25), .CO (n_18));
  ADDFX2 g1219(.A (b[0]), .B (a[0]), .CI (cin), .S (sum[0]), .CO(n_16));
  NAND2BXL g1222(.AN (n_39), .B (n_14), .Y (n_15));
  NAND2BXL g1223(.AN (n_78), .B (n_12), .Y (n_13));
  NAND2BXL g1220(.AN (n_58), .B (n_10), .Y (n_11));
  NAND2BXL g1221(.AN (n_9), .B (n_8), .Y (n_40));
  NAND2BXL g1227(.AN (n_19), .B (n_6), .Y (n_7));
  NAND2BXL g1224(.AN (n_5), .B (n_4), .Y (n_21));
  NAND2BXL g1226(.AN (n_3), .B (n_2), .Y (n_59));
  NAND2BXL g1225(.AN (n_1), .B (n_0), .Y (n_79));
  NAND2XL g1237(.A (b[15]), .B (a[15]), .Y (n_0));
  NAND2XL g1229(.A (b[3]), .B (a[3]), .Y (n_4));
  NOR2XL g1233(.A (a[3]), .B (b[3]), .Y (n_5));
  NAND2XL g1236(.A (b[6]), .B (a[6]), .Y (n_14));
  NAND2XL g1239(.A (b[11]), .B (a[11]), .Y (n_2));
  NOR2XL g1242(.A (a[2]), .B (b[2]), .Y (n_19));
  NOR2XL g1243(.A (a[14]), .B (b[14]), .Y (n_78));
  NOR2XL g1235(.A (a[6]), .B (b[6]), .Y (n_39));
  NAND2XL g1230(.A (b[10]), .B (a[10]), .Y (n_10));
  NOR2XL g1231(.A (a[11]), .B (b[11]), .Y (n_3));
  NAND2XL g1240(.A (b[7]), .B (a[7]), .Y (n_8));
  NOR2XL g1232(.A (a[7]), .B (b[7]), .Y (n_9));
  NAND2XL g1228(.A (b[14]), .B (a[14]), .Y (n_12));
  NOR2XL g1241(.A (a[15]), .B (b[15]), .Y (n_1));
  NAND2XL g1238(.A (b[2]), .B (a[2]), .Y (n_6));
  NOR2XL g1234(.A (a[10]), .B (b[10]), .Y (n_58));
endmodule